module Demodulate(clk, QPSK_out, I_demodulate, Q_demodulate);
  input clk;
  input [9:0] QPSK_out;
  output I_demodulate, Q_demodulate;

endmodule