module adder(clk1, input1, input2, out);
input clk1, input1, input2;
output out;
endmodule